module Debounce(  // edge detect, synchronize to clock, debounce input pushbutton or switch
   input clk, b,  // b is the bouncy pushbutton or switch
   output reg s   // debounced version of pushbutton, synched to clock.
                  // ASSUMES the bouncing continues for less than 2 clock periods  
);

   // insert code here
endmodule